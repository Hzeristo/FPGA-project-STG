module music_3 (
    input clk,
    input rst_n;
    input address,
    output reg[32:0] note
);

//time intervals of each note
localparam              
         
M1=95602,           //1
M11=90253,          //1#
M2=85178,           //2
M21=80386,          //2#
M3=75872,           //3
M4=71633,           //4
M41=67568,          //4#
M5=63775,           //5
M51=60168,          //5#
M6=56818,           //6
M61=53648,          //6#
M7=50607,           //7

H1=47801,           //1
H11=45086,          //1#
H2=42553,           //2
H21=40161,          //2#
H3=37936,           //3
H4=35791,           //4
H41=33784,          //4#
H5=31888,           //5
H51=30102,          //5#
H6=28409,           //6
H61=26810,          //6#
H7=25303,           //7

HH1=23883,
HH2=22543,

D5=127551,          //5
D51=120482,         //5#
D6=113636,          //6
D61=107296,         //6#
D7=101215,          //7
S=2500             //休止符

always @(posedge clk or negedge rst_n) begin
  if (!rst_n) begin
    pre_set <= 0;  
  end else begin
    case(address)
0:pre_set<=M6;
				1:pre_set<=M6;
				2:pre_set<=M2;
				3:pre_set<=M2;
				4:pre_set<=M3;
				5:pre_set<=M3;
				6:pre_set<=D6;
				7:pre_set<=D6;
				8:pre_set<=S;
				9:pre_set<=S;
				10:pre_set<=M6;
				11:pre_set<=M6;
				12:pre_set<=M2;
				13:pre_set<=M2;
				14:pre_set<=M3;
				15:pre_set<=M3;
				16:pre_set<=D6;
				17:pre_set<=D6;
				18:pre_set<=S;
				19:pre_set<=S;
				20:pre_set<=S;
				21:pre_set<=S;
				22:pre_set<=M6;
				23:pre_set<=M6;
				24:pre_set<=M2;
				25:pre_set<=M2;
				26:pre_set<=M3;
				27:pre_set<=M3;
				28:pre_set<=D6;
				29:pre_set<=D6;
				30:pre_set<=S;
				31:pre_set<=S;
				32:pre_set<=M6;
				33:pre_set<=M6;
				34:pre_set<=M2;
				35:pre_set<=M2;
				36:pre_set<=M3;
				37:pre_set<=M3;
				38:pre_set<=D6;
				39:pre_set<=D6;
				40:pre_set<=S;
				41:pre_set<=S;
				42:pre_set<=M6;
				43:pre_set<=M6;
				44:pre_set<=M2;
				45:pre_set<=M2;
				46:pre_set<=M3;
				47:pre_set<=M3;
				48:pre_set<=D6;
				49:pre_set<=D6;
				50:pre_set<=S;
				51:pre_set<=S;
				52:pre_set<=S;
				53:pre_set<=S;
				54:pre_set<=M6;
				55:pre_set<=M6;
				56:pre_set<=M2;
				57:pre_set<=M2;
				58:pre_set<=M3;
				59:pre_set<=M3;
				60:pre_set<=D6;
				61:pre_set<=D6;
				62:pre_set<=S;
				63:pre_set<=S;
				64:pre_set<=M6;
				65:pre_set<=M6;
				66:pre_set<=M2;
				67:pre_set<=M2;
				68:pre_set<=M3;
				69:pre_set<=M3;
				70:pre_set<=D6;
				71:pre_set<=D6;
				72:pre_set<=S;
				73:pre_set<=S;
				74:pre_set<=M6;
				75:pre_set<=M6;
				76:pre_set<=M2;
				77:pre_set<=M2;
				78:pre_set<=M3;
				79:pre_set<=M3;
				80:pre_set<=D6;
				81:pre_set<=D6;
				82:pre_set<=S;
				83:pre_set<=S;
				84:pre_set<=S;
				85:pre_set<=S;
				86:pre_set<=M6;
				87:pre_set<=M6;
				88:pre_set<=M2;
				89:pre_set<=M2;
				90:pre_set<=M3;
				91:pre_set<=M3;
				92:pre_set<=D6;
				93:pre_set<=D6;
				94:pre_set<=S;
				95:pre_set<=S;
				96:pre_set<=M6;
				97:pre_set<=M6;
				98:pre_set<=M2;
				99:pre_set<=M2;
				100:pre_set<=M3;
				101:pre_set<=M3;
				102:pre_set<=D6;
				103:pre_set<=D6;
				104:pre_set<=S;
				105:pre_set<=S;
				106:pre_set<=M6;
				107:pre_set<=M6;
				108:pre_set<=M2;
				109:pre_set<=M2;
				110:pre_set<=M3;
				111:pre_set<=M3;
				112:pre_set<=D6;
				113:pre_set<=D6;
				114:pre_set<=S;
				115:pre_set<=S;
				116:pre_set<=S;
				117:pre_set<=S;
				118:pre_set<=M6;
				119:pre_set<=M6;
				120:pre_set<=M2;
				121:pre_set<=M2;
				122:pre_set<=M3;
				123:pre_set<=M3;
				124:pre_set<=D6;
				125:pre_set<=D6;
				126:pre_set<=S;
				127:pre_set<=S;//主旋律开始
                                128:pre_set<=M3;
				129:pre_set<=M3;
				130:pre_set<=M3;
				131:pre_set<=M3;
				132:pre_set<=M3;
				133:pre_set<=M3;
				134:pre_set<=M3;
				135:pre_set<=M3;
				136:pre_set<=M7;
				137:pre_set<=M7;
				138:pre_set<=M7;
				139:pre_set<=M7;
				140:pre_set<=M7;
				141:pre_set<=M7;
				142:pre_set<=M7;
				143:pre_set<=M7;
				144:pre_set<=H2;
				145:pre_set<=H2;
				146:pre_set<=H2;
				147:pre_set<=H2;
				148:pre_set<=H2;
				149:pre_set<=H2;
				150:pre_set<=H2;
				151:pre_set<=H2;
				152:pre_set<=H1;
				153:pre_set<=H1;
				154:pre_set<=H1;
				155:pre_set<=M7;
				156:pre_set<=M7;
				157:pre_set<=M7;
				158:pre_set<=M5;
				159:pre_set<=M5;
				160:pre_set<=M3;
				161:pre_set<=M3;
				162:pre_set<=M3;
				163:pre_set<=M3;
				164:pre_set<=M3;
				165:pre_set<=M3;
				166:pre_set<=M3;
				167:pre_set<=M3;
				168:pre_set<=M3;
				169:pre_set<=M3;
				170:pre_set<=M3;
				171:pre_set<=M3;
				172:pre_set<=M3;
				173:pre_set<=M3;
				174:pre_set<=M3;
				175:pre_set<=M3;
				176:pre_set<=M3;
				177:pre_set<=M3;
				178:pre_set<=M3;
				179:pre_set<=M3;
				180:pre_set<=M3;
				181:pre_set<=M3;
				182:pre_set<=M3;
				183:pre_set<=M3;
				184:pre_set<=S;
				185:pre_set<=S;
				186:pre_set<=S;
				187:pre_set<=S;
				188:pre_set<=S;
				189:pre_set<=S;
				190:pre_set<=S;
				191:pre_set<=S;
				192:pre_set<=M3;
				193:pre_set<=M3;
				194:pre_set<=M3;
				195:pre_set<=M3;
				196:pre_set<=M3;
				197:pre_set<=M3;
				198:pre_set<=M3;
				199:pre_set<=M3;
				200:pre_set<=M7;
				201:pre_set<=M7;
				202:pre_set<=M7;
				203:pre_set<=M7;
				204:pre_set<=M7;
				205:pre_set<=M7;
				206:pre_set<=M7;
				207:pre_set<=M7;
				208:pre_set<=H2;
				209:pre_set<=H2;
				210:pre_set<=H2;
				211:pre_set<=H2;
				212:pre_set<=H2;
				213:pre_set<=H2;
				214:pre_set<=H2;
				215:pre_set<=H2;
				216:pre_set<=H1;
				217:pre_set<=H1;
				218:pre_set<=H1;
				219:pre_set<=M7;
				220:pre_set<=M7;
				221:pre_set<=M7;
				222:pre_set<=M5;
				223:pre_set<=M5;
				224:pre_set<=M6;
				225:pre_set<=M6;
				226:pre_set<=M6;
				227:pre_set<=M6;
				228:pre_set<=M6;
				229:pre_set<=M6;
				230:pre_set<=M6;
				231:pre_set<=M6;
				232:pre_set<=M6;
				233:pre_set<=M6;
				234:pre_set<=M6;
				235:pre_set<=M6;
				236:pre_set<=M6;
				237:pre_set<=M6;
				238:pre_set<=M6;
				239:pre_set<=M6;
				240:pre_set<=M6;
				241:pre_set<=M6;
				242:pre_set<=M6;
				243:pre_set<=M6;
				244:pre_set<=M6;
				245:pre_set<=M6;
				246:pre_set<=M6;
				247:pre_set<=M6;
				248:pre_set<=S;
				249:pre_set<=S;
				250:pre_set<=S;
				251:pre_set<=S;
				252:pre_set<=S;
				253:pre_set<=S;
				254:pre_set<=S;
				255:pre_set<=S;
				256:pre_set<=H1;
				257:pre_set<=H1;
				258:pre_set<=H1;
				259:pre_set<=H1;
				260:pre_set<=H1;
				261:pre_set<=H1;
				262:pre_set<=H1;
				263:pre_set<=H1;
				264:pre_set<=H2;
				265:pre_set<=H2;
				266:pre_set<=H2;
				267:pre_set<=H2;
				268:pre_set<=H2;
				269:pre_set<=H2;
				270:pre_set<=H2;
				271:pre_set<=H2;
				272:pre_set<=H5;
				273:pre_set<=H5;
				274:pre_set<=H5;
				275:pre_set<=H5;
				276:pre_set<=H5;
				277:pre_set<=H5;
				278:pre_set<=H5;
				279:pre_set<=H5;
				280:pre_set<=H3;
				281:pre_set<=H3;
				282:pre_set<=H3;
				283:pre_set<=H2;
				284:pre_set<=H2;
				285:pre_set<=H2;
				286:pre_set<=M5;
				287:pre_set<=M5;
				288:pre_set<=M6;
				289:pre_set<=M6;
				290:pre_set<=M6;
				291:pre_set<=M6;
				292:pre_set<=M6;
				293:pre_set<=M6;
				294:pre_set<=M6;
				295:pre_set<=M6;
				296:pre_set<=M6;
				297:pre_set<=M6;
				298:pre_set<=M6;
				299:pre_set<=M6;
				300:pre_set<=M6;
				301:pre_set<=M6;
				302:pre_set<=M6;
				303:pre_set<=M6;
				304:pre_set<=S;
				305:pre_set<=S;
				306:pre_set<=S;
				307:pre_set<=S;
				308:pre_set<=S;
				309:pre_set<=S;
				310:pre_set<=S;
				311:pre_set<=S;
				312:pre_set<=H1;
				313:pre_set<=H1;
				314:pre_set<=H1;
				315:pre_set<=H1;
				316:pre_set<=H1;
				317:pre_set<=H1;
				318:pre_set<=H1;
				319:pre_set<=H1;
				320:pre_set<=H5;
				321:pre_set<=H5;
				322:pre_set<=H5;
				323:pre_set<=H5;
				324:pre_set<=H5;
				325:pre_set<=H5;
				326:pre_set<=H5;
				327:pre_set<=H5;
				328:pre_set<=H7;
				329:pre_set<=H7;
				330:pre_set<=H7;
				331:pre_set<=H7;
				332:pre_set<=H7;
				333:pre_set<=H7;
				334:pre_set<=H7;
				335:pre_set<=H7;
				336:pre_set<=HH1;
				337:pre_set<=HH1;
				338:pre_set<=HH1;
				339:pre_set<=H7;
				340:pre_set<=H7;
				341:pre_set<=H7;
				342:pre_set<=H5;
				343:pre_set<=H5;
				344:pre_set<=H6;
				345:pre_set<=H6;
				346:pre_set<=H6;
				347:pre_set<=H6;
				348:pre_set<=H6;
				349:pre_set<=H6;
				350:pre_set<=H6;
				351:pre_set<=H6;
				352:pre_set<=H6;
				353:pre_set<=H6;
				354:pre_set<=H6;
				355:pre_set<=H6;
				356:pre_set<=H6;
				357:pre_set<=H6;
				358:pre_set<=H6;
				359:pre_set<=H6;
				360:pre_set<=M6;
				361:pre_set<=M6;
				362:pre_set<=M6;
				363:pre_set<=M6;
				364:pre_set<=M6;
				365:pre_set<=M6;
				366:pre_set<=M6;
				367:pre_set<=M6;
				368:pre_set<=S;
				369:pre_set<=S;
				370:pre_set<=S;
				371:pre_set<=S;
				372:pre_set<=M3;
				373:pre_set<=M3;
				374:pre_set<=M3;
				375:pre_set<=M3;
				376:pre_set<=D6;
				377:pre_set<=D6;
				378:pre_set<=D6;
				379:pre_set<=D6;
				380:pre_set<=D6;
				381:pre_set<=D6;
				382:pre_set<=D6;
				383:pre_set<=D6;
				384:pre_set<=D6;
				385:pre_set<=D6;
				386:pre_set<=D6;
				387:pre_set<=D6;
				388:pre_set<=D6;
				389:pre_set<=D6;
				390:pre_set<=D6;
				391:pre_set<=D6;
				392:pre_set<=D7;
				393:pre_set<=D7;
				394:pre_set<=D7;
				395:pre_set<=D7;
				396:pre_set<=D7;
				397:pre_set<=D7;
				398:pre_set<=D7;
				399:pre_set<=D7;
				400:pre_set<=D7;
				401:pre_set<=D7;
				402:pre_set<=D7;
				403:pre_set<=D7;
				404:pre_set<=D7;
				405:pre_set<=D7;
				406:pre_set<=D7;
				407:pre_set<=D7;
				408:pre_set<=M1;
				409:pre_set<=M1;
				410:pre_set<=M1;
				411:pre_set<=M1;
				412:pre_set<=M1;
				413:pre_set<=M1;
				414:pre_set<=M1;
				415:pre_set<=M1;
				416:pre_set<=M1;
				417:pre_set<=M1;
				418:pre_set<=M1;
				419:pre_set<=M1;
				420:pre_set<=M1;
				421:pre_set<=M1;
				422:pre_set<=M1;
				423:pre_set<=M1;
				424:pre_set<=M2;
				425:pre_set<=M2;
				426:pre_set<=M2;
				427:pre_set<=M2;
				428:pre_set<=M2;
				429:pre_set<=M2;
				430:pre_set<=M2;
				431:pre_set<=M2;
				432:pre_set<=M3;
				433:pre_set<=M3;
				434:pre_set<=M3;
				435:pre_set<=M3;
				436:pre_set<=M5;
				437:pre_set<=M5;
				438:pre_set<=M5;
				439:pre_set<=M5;
				440:pre_set<=M6;
				441:pre_set<=M6;
				442:pre_set<=M6;
				443:pre_set<=M6;
				444:pre_set<=M6;
				445:pre_set<=M6;
				446:pre_set<=M6;
				447:pre_set<=M6;
				448:pre_set<=M5;
				449:pre_set<=M5;
				450:pre_set<=M5;
				451:pre_set<=M5;
				452:pre_set<=M6;
				453:pre_set<=M6;
				454:pre_set<=M6;
				455:pre_set<=M6;
				456:pre_set<=H1;
				457:pre_set<=H1;
				458:pre_set<=H1;
				459:pre_set<=H1;
				460:pre_set<=M7;
				461:pre_set<=M7;
				462:pre_set<=M7;
				463:pre_set<=M7;
				464:pre_set<=M2;
				465:pre_set<=M2;
				466:pre_set<=M2;
				467:pre_set<=M2;
				468:pre_set<=M5;
				469:pre_set<=M5;
				470:pre_set<=M5;
				471:pre_set<=M5;
				472:pre_set<=M3;
				473:pre_set<=M3;
				474:pre_set<=M3;
				475:pre_set<=M3;
				476:pre_set<=M3;
				477:pre_set<=M3;
				478:pre_set<=M3;
				479:pre_set<=M3;
				480:pre_set<=M3;
				481:pre_set<=M3;
				482:pre_set<=M3;
				483:pre_set<=M3;
				484:pre_set<=M3;
				485:pre_set<=M3;
				486:pre_set<=M3;
				487:pre_set<=M3;
				488:pre_set<=M3;
				489:pre_set<=M3;
				490:pre_set<=M3;
				491:pre_set<=M3;
				492:pre_set<=M3;
				493:pre_set<=M3;
				494:pre_set<=S;
				495:pre_set<=S;
				496:pre_set<=M3;
				497:pre_set<=M3;
				498:pre_set<=M3;
				499:pre_set<=M3;
				500:pre_set<=M3;
				501:pre_set<=M3;
				502:pre_set<=M3;
				503:pre_set<=M3;
				504:pre_set<=D6;
				505:pre_set<=D6;
				506:pre_set<=D6;
				507:pre_set<=D6;
				508:pre_set<=D6;
				509:pre_set<=D6;
				510:pre_set<=D6;
				511:pre_set<=D6;
				512:pre_set<=D6;
				513:pre_set<=D6;
				514:pre_set<=D6;
				515:pre_set<=D6;
				516:pre_set<=D6;
				517:pre_set<=D6;
				518:pre_set<=D6;
				519:pre_set<=D6;
				520:pre_set<=D7;
				521:pre_set<=D7;
				522:pre_set<=D7;
				523:pre_set<=D7;
				524:pre_set<=D7;
				525:pre_set<=D7;
				526:pre_set<=D7;
				527:pre_set<=D7;
				528:pre_set<=D7;
				529:pre_set<=D7;
				530:pre_set<=D7;
				531:pre_set<=D7;
				532:pre_set<=D7;
				533:pre_set<=D7;
				534:pre_set<=D7;
				535:pre_set<=D7;
				536:pre_set<=M1;
				537:pre_set<=M1;
				538:pre_set<=M1;
				539:pre_set<=M1;
				540:pre_set<=M1;
				541:pre_set<=M1;
				542:pre_set<=M1;
				543:pre_set<=M1;
				544:pre_set<=M1;
				545:pre_set<=M1;
				546:pre_set<=M1;
				547:pre_set<=M1;
				548:pre_set<=M1;
				549:pre_set<=M1;
				550:pre_set<=M1;
				551:pre_set<=M1;
				552:pre_set<=M2;
				553:pre_set<=M2;
				554:pre_set<=M2;
				555:pre_set<=M2;
				556:pre_set<=M2;
				557:pre_set<=M2;
				558:pre_set<=M2;
				559:pre_set<=M2;
				560:pre_set<=M3;
				561:pre_set<=M3;
				562:pre_set<=M3;
				563:pre_set<=M3;
				564:pre_set<=M5;
				565:pre_set<=M5;
				566:pre_set<=M5;
				567:pre_set<=M5;
				568:pre_set<=M6;
				569:pre_set<=M6;
				570:pre_set<=M6;
				571:pre_set<=M6;
				572:pre_set<=M6;
				573:pre_set<=M6;
				574:pre_set<=M6;
				575:pre_set<=M6;
				576:pre_set<=M5;
				577:pre_set<=M5;
				578:pre_set<=M5;
				579:pre_set<=M5;
				580:pre_set<=M6;
				581:pre_set<=M6;
				582:pre_set<=M6;
				583:pre_set<=M6;
				584:pre_set<=H1;
				585:pre_set<=H1;
				586:pre_set<=H1;
				587:pre_set<=H1;
				588:pre_set<=M7;
				589:pre_set<=M7;
				590:pre_set<=M7;
				591:pre_set<=M7;
				592:pre_set<=M5;
				593:pre_set<=M5;
				594:pre_set<=M5;
				595:pre_set<=M5;
				596:pre_set<=M5;
				597:pre_set<=M5;
				598:pre_set<=M5;
				599:pre_set<=M5;
				600:pre_set<=M6;
				601:pre_set<=M6;
				602:pre_set<=M6;
				603:pre_set<=M6;
				604:pre_set<=M6;
				605:pre_set<=M6;
				606:pre_set<=M6;
				607:pre_set<=M6;
				608:pre_set<=M6;
				609:pre_set<=M6;
				610:pre_set<=M6;
				611:pre_set<=M6;
				612:pre_set<=M6;
				613:pre_set<=M6;
				614:pre_set<=M6;
				615:pre_set<=M6;
				616:pre_set<=M6;
				617:pre_set<=M6;
				618:pre_set<=M6;
				619:pre_set<=M6;
				620:pre_set<=M6;
				621:pre_set<=M6;
				622:pre_set<=M6;
				623:pre_set<=M6;
				624:pre_set<=S;
				625:pre_set<=S;
				626:pre_set<=S;
				627:pre_set<=S;
				628:pre_set<=S;
				629:pre_set<=S;
				630:pre_set<=S;
				631:pre_set<=S;
				632:pre_set<=D6;
				633:pre_set<=D6;
				634:pre_set<=D6;
				635:pre_set<=D6;
				636:pre_set<=D6;
				637:pre_set<=D6;
				638:pre_set<=D6;
				639:pre_set<=D6;
				640:pre_set<=D6;
				641:pre_set<=D6;
				642:pre_set<=D6;
				643:pre_set<=D6;
				644:pre_set<=D6;
				645:pre_set<=D6;
				646:pre_set<=D6;
				647:pre_set<=D6;
				648:pre_set<=D7;
				649:pre_set<=D7;
				650:pre_set<=D7;
				651:pre_set<=D7;
				652:pre_set<=D7;
				653:pre_set<=D7;
				654:pre_set<=D7;
				655:pre_set<=D7;
				656:pre_set<=D7;
				657:pre_set<=D7;
				658:pre_set<=D7;
				659:pre_set<=D7;
				660:pre_set<=D7;
				661:pre_set<=D7;
				662:pre_set<=D7;
				663:pre_set<=D7;
				664:pre_set<=M1;
				665:pre_set<=M1;
				666:pre_set<=M1;
				667:pre_set<=M1;
				668:pre_set<=M1;
				669:pre_set<=M1;
				670:pre_set<=M1;
				671:pre_set<=M1;
				672:pre_set<=M1;
				673:pre_set<=M1;
				674:pre_set<=M1;
				675:pre_set<=M1;
				676:pre_set<=M1;
				677:pre_set<=M1;
				678:pre_set<=M1;
				679:pre_set<=M1;
				680:pre_set<=M2;
				681:pre_set<=M2;
				682:pre_set<=M2;
				683:pre_set<=M2;
				684:pre_set<=M2;
				685:pre_set<=M2;
				686:pre_set<=M2;
				687:pre_set<=M2;
				688:pre_set<=M3;
				689:pre_set<=M3;
				690:pre_set<=M3;
				691:pre_set<=M3;
				692:pre_set<=M5;
				693:pre_set<=M5;
				694:pre_set<=M5;
				695:pre_set<=M5;
				696:pre_set<=M6;
				697:pre_set<=M6;
				698:pre_set<=M6;
				699:pre_set<=M6;
				700:pre_set<=M6;
				701:pre_set<=M6;
				702:pre_set<=M6;
				703:pre_set<=M6;
				704:pre_set<=M5;
				705:pre_set<=M5;
				706:pre_set<=M5;
				707:pre_set<=M5;
				708:pre_set<=M6;
				709:pre_set<=M6;
				710:pre_set<=M6;
				711:pre_set<=M6;
				712:pre_set<=H1;
				713:pre_set<=H1;
				714:pre_set<=H1;
				715:pre_set<=H1;
				716:pre_set<=M7;
				717:pre_set<=M7;
				718:pre_set<=M7;
				719:pre_set<=M7;
				720:pre_set<=M2;
				721:pre_set<=M2;
				722:pre_set<=M2;
				723:pre_set<=M2;
				724:pre_set<=M5;
				725:pre_set<=M5;
				726:pre_set<=M5;
				727:pre_set<=M5;
				728:pre_set<=M3;
				729:pre_set<=M3;
				730:pre_set<=M3;
				731:pre_set<=M3;
				732:pre_set<=M3;
				733:pre_set<=M3;
				734:pre_set<=M3;
				735:pre_set<=M3;
				736:pre_set<=M3;
				737:pre_set<=M3;
				738:pre_set<=M3;
				739:pre_set<=M3;
				740:pre_set<=M3;
				741:pre_set<=M3;
				742:pre_set<=M3;
				743:pre_set<=M3;
				744:pre_set<=M3;
				745:pre_set<=M3;
				746:pre_set<=M3;
				747:pre_set<=M3;
				748:pre_set<=M3;
				749:pre_set<=M3;
				750:pre_set<=S;
				751:pre_set<=S;
				752:pre_set<=M3;
				753:pre_set<=M3;
				754:pre_set<=M3;
				755:pre_set<=M3;
				756:pre_set<=M3;
				757:pre_set<=M3;
				758:pre_set<=M3;
				759:pre_set<=M3;
				760:pre_set<=D6;
				761:pre_set<=D6;
				762:pre_set<=D6;
				763:pre_set<=D6;
				764:pre_set<=D6;
				765:pre_set<=D6;
				766:pre_set<=D6;
				767:pre_set<=D6;
				768:pre_set<=D6;
				769:pre_set<=D6;
				770:pre_set<=D6;
				771:pre_set<=D6;
				772:pre_set<=D6;
				773:pre_set<=D6;
				774:pre_set<=D6;
				775:pre_set<=D6;
				776:pre_set<=D7;
				777:pre_set<=D7;
				778:pre_set<=D7;
				779:pre_set<=D7;
				780:pre_set<=D7;
				781:pre_set<=D7;
				782:pre_set<=D7;
				783:pre_set<=D7;
				784:pre_set<=D7;
				785:pre_set<=D7;
				786:pre_set<=D7;
				787:pre_set<=D7;
				788:pre_set<=D7;
				789:pre_set<=D7;
				790:pre_set<=D7;
				791:pre_set<=D7;
				792:pre_set<=M1;
				793:pre_set<=M1;
				794:pre_set<=M1;
				795:pre_set<=M1;
				796:pre_set<=M1;
				797:pre_set<=M1;
				798:pre_set<=M1;
				799:pre_set<=M1;
				800:pre_set<=M1;
				801:pre_set<=M1;
				802:pre_set<=M1;
				803:pre_set<=M1;
				804:pre_set<=M1;
				805:pre_set<=M1;
				806:pre_set<=M1;
				807:pre_set<=M1;
				808:pre_set<=M2;
				809:pre_set<=M2;
				810:pre_set<=M2;
				811:pre_set<=M2;
				812:pre_set<=M2;
				813:pre_set<=M2;
				814:pre_set<=M2;
				815:pre_set<=M2;
				816:pre_set<=M3;
				817:pre_set<=M3;
				818:pre_set<=M3;
				819:pre_set<=M3;
				820:pre_set<=M5;
				821:pre_set<=M5;
				822:pre_set<=M5;
				823:pre_set<=M5;
				824:pre_set<=M6;
				825:pre_set<=M6;
				826:pre_set<=M6;
				827:pre_set<=M6;
				828:pre_set<=M6;
				829:pre_set<=M6;
				830:pre_set<=M6;
				831:pre_set<=M6;
				832:pre_set<=M5;
				833:pre_set<=M5;
				834:pre_set<=M5;
				835:pre_set<=M5;
				836:pre_set<=M6;
				837:pre_set<=M6;
				838:pre_set<=M6;
				839:pre_set<=M6;
				840:pre_set<=H1;
				841:pre_set<=H1;
				842:pre_set<=H1;
				843:pre_set<=H1;
				844:pre_set<=M7;
				845:pre_set<=M7;
				846:pre_set<=M7;
				847:pre_set<=M7;
				848:pre_set<=M5;
				849:pre_set<=M5;
				850:pre_set<=M5;
				851:pre_set<=M5;
				852:pre_set<=M5;
				853:pre_set<=M5;
				854:pre_set<=M5;
				855:pre_set<=M5;
				856:pre_set<=M6;
				857:pre_set<=M6;
				858:pre_set<=M6;
				859:pre_set<=M6;
				860:pre_set<=M6;
				861:pre_set<=M6;
				862:pre_set<=M6;
				863:pre_set<=M6;
				864:pre_set<=M6;
				865:pre_set<=M6;
				866:pre_set<=M6;
				867:pre_set<=M6;
				868:pre_set<=M6;
				869:pre_set<=M6;
				870:pre_set<=M6;
				871:pre_set<=M6;
				872:pre_set<=M6;
				873:pre_set<=M6;
				874:pre_set<=M6;
				875:pre_set<=M6;
				876:pre_set<=M6;
				877:pre_set<=M6;
				878:pre_set<=M6;
				879:pre_set<=M6;
				880:pre_set<=S;
				881:pre_set<=S;
				882:pre_set<=S;
				883:pre_set<=S;
				884:pre_set<=S;
				885:pre_set<=S;
				886:pre_set<=S;
				887:pre_set<=S;//主旋律结束
				888:pre_set<=M6;
				889:pre_set<=M6;
				890:pre_set<=S;
				891:pre_set<=S;
				892:pre_set<=S;
				893:pre_set<=S;
				894:pre_set<=M7;
				895:pre_set<=H1;
				896:pre_set<=H2;
				897:pre_set<=H2;
				898:pre_set<=H3;
				899:pre_set<=H3;
				900:pre_set<=M6;
				901:pre_set<=M6;
				902:pre_set<=M6;
				903:pre_set<=M6;
				904:pre_set<=M3;
				905:pre_set<=M3;
				906:pre_set<=S;
				907:pre_set<=S;
				908:pre_set<=S;
				909:pre_set<=S;
				910:pre_set<=M4;
				911:pre_set<=M5;
				912:pre_set<=M6;
				913:pre_set<=M6;
				914:pre_set<=M7;
				915:pre_set<=M7;
				916:pre_set<=M3;
				917:pre_set<=M3;
				918:pre_set<=M3;
				919:pre_set<=M3;
				920:pre_set<=M4;
				921:pre_set<=M4;
				922:pre_set<=M5;
				923:pre_set<=M5;
				924:pre_set<=M6;
				925:pre_set<=M6;
				926:pre_set<=M3;
				927:pre_set<=M4;
				928:pre_set<=M5;
				929:pre_set<=M5;
				930:pre_set<=M6;
				931:pre_set<=M6;
				932:pre_set<=M7;
				933:pre_set<=M7;
				934:pre_set<=M5;
				935:pre_set<=M5;
				936:pre_set<=H1;
				937:pre_set<=H1;
				938:pre_set<=M7;
				939:pre_set<=M7;
				940:pre_set<=M5;
				941:pre_set<=M5;
				942:pre_set<=M6;
				943:pre_set<=M6;
				944:pre_set<=M3;
				945:pre_set<=M3;
				946:pre_set<=M5;
				947:pre_set<=M5;
				948:pre_set<=M2;
				949:pre_set<=M2;
				950:pre_set<=M2;
				951:pre_set<=M2;
				952:pre_set<=M6;
				953:pre_set<=M6;
				954:pre_set<=S;
				955:pre_set<=S;
				956:pre_set<=S;
				957:pre_set<=S;
				958:pre_set<=M7;
				959:pre_set<=H1;
				960:pre_set<=H2;
				961:pre_set<=H2;
				962:pre_set<=H3;
				963:pre_set<=H3;
				964:pre_set<=M6;
				965:pre_set<=M6;
				966:pre_set<=M6;
				967:pre_set<=M6;
				968:pre_set<=M3;
				969:pre_set<=M3;
				970:pre_set<=S;
				971:pre_set<=S;
				972:pre_set<=S;
				973:pre_set<=S;
				974:pre_set<=M4;
				975:pre_set<=M5;
				976:pre_set<=M6;
				977:pre_set<=M6;
				978:pre_set<=M7;
				979:pre_set<=M7;
				980:pre_set<=M3;
				981:pre_set<=M3;
				982:pre_set<=M3;
				983:pre_set<=M3;
				984:pre_set<=M4;
				985:pre_set<=M4;
				986:pre_set<=M5;
				987:pre_set<=M5;
				988:pre_set<=M6;
				989:pre_set<=M6;
				990:pre_set<=M3;
				991:pre_set<=M3;
				992:pre_set<=H1;
				993:pre_set<=H1;
				994:pre_set<=M7;
				995:pre_set<=M7;
				996:pre_set<=M5;
				997:pre_set<=M5;
				998:pre_set<=M6;
				999:pre_set<=M6;
				1000:pre_set<=M51;
				1001:pre_set<=M51;
				1002:pre_set<=M51;
				1003:pre_set<=M5;
				1004:pre_set<=M5;
				1005:pre_set<=S;
				1006:pre_set<=M5;
				1007:pre_set<=M6;
				1008:pre_set<=M7;
				1009:pre_set<=M7;
				1010:pre_set<=M7;
				1011:pre_set<=M7;
				1012:pre_set<=M7;
				1013:pre_set<=M7;
				1014:pre_set<=M7;
				1015:pre_set<=M7;
				1016:pre_set<=M6;
				1017:pre_set<=M6;
				1018:pre_set<=S;
				1019:pre_set<=S;
				1020:pre_set<=S;
				1021:pre_set<=S;
				1022:pre_set<=M7;
				1023:pre_set<=H1;
				default:pre_set<=0;
    endcase
  end
end

endmodule