module music_2 (
    input clk,
    input rst_n;
    input address,
    output reg[32:0] note
);

//time intervals of each note
localparam              
            M1=95602,           //1
            M11=90253,          //1#
	        M2=85178,           //2
		    M21=80386,         //2#
	        M3=75872,           //3
	        M4=71633,           //4
		    M41=67568,          //4#
	        M5=63775,           //5
	    	M51=60168,          //5#
    	    M6=56818,           //6
		    M61=53648,          //6#
	        M7=50607,           //7
      //high key
			H1=47801,           //1
			H11=45086,           //1#
			H2=42553,           //2
			H21=40161,           //2#
			H3=37936,           //3
			H4=35791,           //4
			H41=33784,           //4#
			H5=31888,           //5
			H51=30102,           //5#
			H6=28409,          //6
			H61=26810,          //6#
			H7=25303,          //7

			//更高音
	        HH1=23883,
	        HH2=22543,

			//low key
			D5=127551,          //5
			D51=120482,         //5#
			D6=113636,          //6
			D61=107296,         //6#
			D7=101215,          //7
			S=2500;             //休止符


always @(posedge clk or negedge rst_n) begin
  if (!rst_n) begin
    pre_set <= 0;  
  end else begin
    case(address)
                0:pre_set<=M6;
				1:pre_set<=M6;
				2:pre_set<=M1;
				3:pre_set<=M6;
				4:pre_set<=M1;
				5:pre_set<=M1;
				6:pre_set<=M6;
				7:pre_set<=S;
				8:pre_set<=M6;
				9:pre_set<=M6;
				10:pre_set<=M1;
				11:pre_set<=M6;
				12:pre_set<=M1;
				13:pre_set<=M1;
				14:pre_set<=M6;
				15:pre_set<=M6;
				16:pre_set<=D7;
				17:pre_set<=D7;
				18:pre_set<=M5;
				19:pre_set<=M5;
				20:pre_set<=M2;
				21:pre_set<=M2;
				22:pre_set<=M7;
				23:pre_set<=M7;
				24:pre_set<=M6;
				25:pre_set<=M6;
				26:pre_set<=M1;
				27:pre_set<=M6;
				28:pre_set<=M1;
				29:pre_set<=M1;
				30:pre_set<=M6;
				31:pre_set<=S;
				32:pre_set<=M6;
				33:pre_set<=M6;
				34:pre_set<=M1;
				35:pre_set<=M6;
				36:pre_set<=M1;
				37:pre_set<=M1;
				38:pre_set<=M6;
				39:pre_set<=S;
				40:pre_set<=M6;
				41:pre_set<=M6;
				42:pre_set<=M1;
				43:pre_set<=M6;
				44:pre_set<=M1;
				45:pre_set<=M1;
				46:pre_set<=M6;
				47:pre_set<=M6;
				48:pre_set<=D7;
				49:pre_set<=D7;
				50:pre_set<=M5;
				51:pre_set<=M5;
				52:pre_set<=M2;
				53:pre_set<=M2;
				54:pre_set<=M7;
				55:pre_set<=M7;
				56:pre_set<=H1;
				57:pre_set<=H1;
				58:pre_set<=M3;
				59:pre_set<=H1;
				60:pre_set<=M3;
				61:pre_set<=M3;
				62:pre_set<=H1;
				63:pre_set<=H1;
				64:pre_set<=M6;
				65:pre_set<=M6;
				66:pre_set<=M1;
				67:pre_set<=M6;
				68:pre_set<=M1;
				69:pre_set<=M1;
				70:pre_set<=M6;
				71:pre_set<=S;
				72:pre_set<=M6;
				73:pre_set<=M6;
				74:pre_set<=M1;
				75:pre_set<=M6;
				76:pre_set<=M1;
				77:pre_set<=M1;
				78:pre_set<=M6;
				79:pre_set<=M6;
				80:pre_set<=D7;
				81:pre_set<=D7;
				82:pre_set<=M5;
				83:pre_set<=M5;
				84:pre_set<=M2;
				85:pre_set<=M2;
				86:pre_set<=M7;
				87:pre_set<=M7;
				88:pre_set<=M51;
				89:pre_set<=M51;
				90:pre_set<=D7;
				91:pre_set<=M51;
				92:pre_set<=D7;
				93:pre_set<=D7;
				94:pre_set<=M51;
				95:pre_set<=M51;
				96:pre_set<=M6;
				97:pre_set<=M6;
				98:pre_set<=M1;
				99:pre_set<=M6;
				100:pre_set<=M1;
				101:pre_set<=M1;
				102:pre_set<=M6;
				103:pre_set<=S;
				104:pre_set<=M6;
				105:pre_set<=M6;
				106:pre_set<=M1;
				107:pre_set<=M6;
				108:pre_set<=M1;
				109:pre_set<=M1;
				110:pre_set<=M6;
				111:pre_set<=M6;
				112:pre_set<=D7;
				113:pre_set<=D7;
				114:pre_set<=M5;
				115:pre_set<=M5;
				116:pre_set<=M2;
				117:pre_set<=M2;
				118:pre_set<=M7;
				119:pre_set<=M7;
				120:pre_set<=M51;
				121:pre_set<=M51;
				122:pre_set<=D61;
				123:pre_set<=D61;
				124:pre_set<=M1;//主旋律开始
				125:pre_set<=M1;
				126:pre_set<=M21;
				127:pre_set<=M21;
                128:pre_set<=H2;
				129:pre_set<=H2;
				130:pre_set<=H2;
				131:pre_set<=H2;
				132:pre_set<=H2;
				133:pre_set<=H2;
				134:pre_set<=H3;
				135:pre_set<=H3;
				136:pre_set<=H2;
				137:pre_set<=H2;
				138:pre_set<=H3;
				139:pre_set<=H3;
				140:pre_set<=H5;
				141:pre_set<=H5;
				142:pre_set<=H3;
				143:pre_set<=H3;
				144:pre_set<=H2;
				145:pre_set<=H2;
				146:pre_set<=H3;
				147:pre_set<=H3;
				148:pre_set<=M6;
				149:pre_set<=M6;
				150:pre_set<=M6;
				151:pre_set<=M6;
				152:pre_set<=S;
				153:pre_set<=S;
				154:pre_set<=M5;
				155:pre_set<=M5;
				156:pre_set<=M6;
				157:pre_set<=M6;
				158:pre_set<=H1;
				159:pre_set<=H1;
				160:pre_set<=H2;
				161:pre_set<=H2;
				162:pre_set<=H2;
				163:pre_set<=H2;
				164:pre_set<=H2;
				165:pre_set<=H2;
				166:pre_set<=H3;
				167:pre_set<=H3;
				168:pre_set<=H5;
				169:pre_set<=H5;
				170:pre_set<=H3;
				171:pre_set<=H3;
				172:pre_set<=H2;
				173:pre_set<=H2;
				174:pre_set<=H3;
				175:pre_set<=H3;
				176:pre_set<=H6;
				177:pre_set<=H6;
				178:pre_set<=H6;
				179:pre_set<=H6;
				180:pre_set<=H6;
				181:pre_set<=H6;
				182:pre_set<=H6;
				183:pre_set<=H6;
				184:pre_set<=S;
				185:pre_set<=S;
				186:pre_set<=H3;
				187:pre_set<=H3;
				188:pre_set<=H6;
				189:pre_set<=H6;
				190:pre_set<=H7;
				191:pre_set<=H7;
				192:pre_set<=HH1;
				193:pre_set<=HH1;
				194:pre_set<=HH1;
				195:pre_set<=HH1;
				196:pre_set<=HH1;
				197:pre_set<=HH1;
				198:pre_set<=HH2;//未定义
				199:pre_set<=HH2;
				200:pre_set<=H7;
				201:pre_set<=H7;
				202:pre_set<=HH1;
				203:pre_set<=HH1;
				204:pre_set<=H7;
				205:pre_set<=H7;
				206:pre_set<=H5;
				207:pre_set<=H5;
				208:pre_set<=H2;
				209:pre_set<=H2;
				210:pre_set<=H3;
				211:pre_set<=H3;
				212:pre_set<=M6;
				213:pre_set<=M6;
				214:pre_set<=M6;
				215:pre_set<=M6;
				216:pre_set<=S;
				217:pre_set<=S;
				218:pre_set<=M3;
				219:pre_set<=M3;
				220:pre_set<=M6;
				221:pre_set<=M6;
				222:pre_set<=M7;
				223:pre_set<=M7;
				224:pre_set<=H1;
				225:pre_set<=H1;
				226:pre_set<=H1;
				227:pre_set<=H1;
				228:pre_set<=H1;
				229:pre_set<=H1;
				230:pre_set<=H3;
				231:pre_set<=H3;
				232:pre_set<=H2;
				233:pre_set<=H2;
				234:pre_set<=H1;
				235:pre_set<=H1;
				236:pre_set<=M7;
				237:pre_set<=M7;
				238:pre_set<=M7;
				239:pre_set<=M7;
				240:pre_set<=M6;
				241:pre_set<=M6;
				242:pre_set<=M6;
				243:pre_set<=M6;
				244:pre_set<=M6;
				245:pre_set<=M6;
				246:pre_set<=M6;
				247:pre_set<=M6;
				248:pre_set<=S;
				249:pre_set<=S;
				250:pre_set<=M5;
				251:pre_set<=M5;
				252:pre_set<=M6;
				253:pre_set<=M6;
				254:pre_set<=H1;
				255:pre_set<=H1;
				256:pre_set<=H2;
				257:pre_set<=H2;
				258:pre_set<=H2;
				259:pre_set<=H2;
				260:pre_set<=H2;
				261:pre_set<=H2;
				262:pre_set<=H3;
				263:pre_set<=H3;
				264:pre_set<=H2;
				265:pre_set<=H2;
				266:pre_set<=H3;
				267:pre_set<=H3;
				268:pre_set<=H5;
				269:pre_set<=H5;
				270:pre_set<=H3;
				271:pre_set<=H3;
				272:pre_set<=H2;
				273:pre_set<=H2;
				274:pre_set<=H3;
				275:pre_set<=H3;
				276:pre_set<=M6;
				277:pre_set<=M6;
				278:pre_set<=M6;
				279:pre_set<=M6;
				280:pre_set<=S;
				281:pre_set<=S;
				282:pre_set<=M5;
				283:pre_set<=M5;
				284:pre_set<=M6;
				285:pre_set<=M6;
				286:pre_set<=H1;
				287:pre_set<=H1;
				288:pre_set<=H2;
				289:pre_set<=H2;
				290:pre_set<=H2;
				291:pre_set<=H2;
				292:pre_set<=H2;
				293:pre_set<=H2;
				294:pre_set<=H3;
				295:pre_set<=H3;
				296:pre_set<=H5;
				297:pre_set<=H5;
				298:pre_set<=H3;
				299:pre_set<=H3;
				300:pre_set<=H2;
				301:pre_set<=H2;
				302:pre_set<=H3;
				303:pre_set<=H3;
				304:pre_set<=H6;
				305:pre_set<=H6;
				306:pre_set<=H6;
				307:pre_set<=H6;
				308:pre_set<=H6;
				309:pre_set<=H6;
				310:pre_set<=H6;
				311:pre_set<=H6;
				312:pre_set<=S;
				313:pre_set<=S;
				314:pre_set<=H3;
				315:pre_set<=H3;
				316:pre_set<=H6;
				317:pre_set<=H6;
				318:pre_set<=H7;
				319:pre_set<=H7;
				320:pre_set<=HH1;
				321:pre_set<=HH1;
				322:pre_set<=HH1;
				323:pre_set<=HH1;
				324:pre_set<=HH1;
				325:pre_set<=HH1;
				326:pre_set<=HH2;
				327:pre_set<=HH2;
				328:pre_set<=H7;
				329:pre_set<=H7;
				330:pre_set<=HH1;
				331:pre_set<=HH1;
				332:pre_set<=H7;
				333:pre_set<=H7;
				334:pre_set<=H5;
				335:pre_set<=H5;
				336:pre_set<=H2;
				337:pre_set<=H2;
				338:pre_set<=H3;
				339:pre_set<=H3;
				340:pre_set<=M6;
				341:pre_set<=M6;
				342:pre_set<=M6;
				343:pre_set<=M6;
				344:pre_set<=S;
				345:pre_set<=S;
				346:pre_set<=M3;
				347:pre_set<=M3;
				348:pre_set<=M6;
				349:pre_set<=M6;
				350:pre_set<=M7;
				351:pre_set<=M7;
				352:pre_set<=H1;
				353:pre_set<=H1;
				354:pre_set<=H1;
				355:pre_set<=H1;
				356:pre_set<=H1;
				357:pre_set<=H1;
				358:pre_set<=H3;
				359:pre_set<=H3;
				360:pre_set<=H2;
				361:pre_set<=H2;
				362:pre_set<=H1;
				363:pre_set<=H1;
				364:pre_set<=M7;
				365:pre_set<=M7;
				366:pre_set<=M7;
				367:pre_set<=M7;
				368:pre_set<=M6;
				369:pre_set<=M6;
				370:pre_set<=M6;
				371:pre_set<=M6;
				372:pre_set<=M6;
				373:pre_set<=M6;
				374:pre_set<=M6;
				375:pre_set<=M6;//finish
				376:pre_set<=M6;
				377:pre_set<=M6;
				378:pre_set<=S;
				379:pre_set<=S;
				380:pre_set<=S;
				381:pre_set<=S;
				382:pre_set<=S;
				383:pre_set<=S;
				default:pre_set<=0;
    endcase
  end
end

endmodule